component traffic_light.CDiagMessage

endpoints {
    message : traffic_light.IDiagMessage
}