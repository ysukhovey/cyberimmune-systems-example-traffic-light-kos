component traffic_light.CCode

endpoints {
    mode : traffic_light.ICode
}
