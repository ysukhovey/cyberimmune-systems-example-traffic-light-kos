component traffic_light.CCode

endpoints {
    code : traffic_light.ICode
}
