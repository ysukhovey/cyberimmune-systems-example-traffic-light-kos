/* Definition of the `Mode` component. */

component traffic_light.CMode

endpoints {
    /* Declaration of a named implementation of the "Mode" interface. */
    mode : traffic_light.IMode
}
